module barrier_data (
	input [7:0] cnt,
	
	output reg [2:0] barrier_out
);

always @ (*) begin
	case (cnt)
		0,1,2,3,4,5,6,7,8,9:
			barrier_out <= 3'b000;
		24,96,156,135,196,4586,1316,16656,13561,5846,156,31,65,349,13,113,519,1323,2189,6351,3613,1513:
			barrier_out <= 3'b110;
		35,99,13,416,151,6156,84,151456,123,561,156,541,31,616,115,325,1616,1565,51,1066,3226,1321,6156,515,361,333,156498,56496,1415,31165,3113,2613,4488,8998,1156,1316,684,4651,35,64,61,43,134,869,183,93,846,4614,463,123,66,464898,4654,1653,1468,46,146,311,638,719,813,5113,446,94,464,54614,98,121,368,461,3615,49,56,613,7564,961,1583,933,413,391,411,6115,113,987,156,9113,774,748,491,1345,3648,871:
			barrier_out <= 3'b010;
		118,928,436,411,561,32,61,612,121,321,133,815,5661,95,561,6132,273,312,561,498,79,444,918,268,614,4011,1126,163,1635,50980,194,319,10484,159,1662,1015,406,480,29,601,80,1156,2104,485,350,486,3690,1406,8060,1305,1056,151,102,16,266,321,610,151,32312,630,36,13,10,5610,9010,305,156,1568,801,46,706,71,681,756:
			barrier_out <= 3'b100;
		12,563,35,665,784,81,87,44,9646,555,54546,113,66,849,471,123,346,16,48,146,511,654,658,131,464,649,414196,879,478,641,99,41,49,14,1916,46,849,481,63105,196,561,4806,561,3058,620,90,06,610,641,676,689,498,96:
			barrier_out <= 3'b001;
		60:
			barrier_out <= 3'b011;
		24:
			barrier_out <= 3'b101;

		default:
			barrier_out <= 3'b000;
	endcase
end

endmodule
